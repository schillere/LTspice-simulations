PID1.CIR - PID CONTROLLER
*
* SET POINT
VSET	1	0	PWL(0MS 0MV   1MS 10V   2000MS 10V)
RSET	1	0	1MEG
*
* CALCULATE ERROR
EERROR	2 0	1 12	1
RERROR	2	0	1MEG
*
* P - PROPORTIONAL TERM
EP	3 0	2 0 1
RP	3	0	1MEG
*
* I - INTEGRAL TERM
GI	0 4	2 0 1
C1	4	0	1
R1	4	0	1MEG
*
* D - DERIVATIVE TERM
GD	0 5	2 0 1
L1	5	0	1
*
* ADD PID TERMS, ADJUST PID MULTIPLIERS
EPID	6 0	POLY(3) (3,0) (4,0) (5,0) 0 1 0 0
*EPID	6 0	VALUE = { 1*V(3) + 0*V(4) + 0*V(5) }
RPID	6	0	1MEG
*
* AMPLIFIER
EAMP	7 0	6 0	1
RAMP	7	0	1MEG
*
* PROCESS BLOCK WITH TIME LAG (PHASE SHIFT)
EOUT	8 0	7 0	100
RP1	8	9	100K
CP1	9	0	1UF
RP2	9	10	100K
CP2	10	0	1UF
*
* SENSOR BLOCK WITH TIME LAG
ESENSOR	11 0	10 0	0.01
RP3	11	12	10K
CP3	12	0	1UF
*
* ANALYSIS
.TRAN 	10MS 2000MS
*
* VIEW RESULTS
*.PRINT TRAN	V(1) V(12)
.PROBE
.END

DC_MOTOR_MODEL.CIR
*
V_AMP	1	0	AC	1 	PWL(0MS 0 50MS 0 50.1MS 10 150MS 10 150.1MS 0)
*
* MOTOR VOLTAGE
RA	1	2	0.5
LA	2	3	0.0015
H_EMF	3 4	VSENSE2	0.05
VSENSE1	4	0	DC 0V
*
* MOTOR TORQUE BASED ON INERTIA AND FRICTION
H_TORQ	6 0	VSENSE1	0.05
LJ	6	7	0.00025
RB	7	8	0.0001
VSENSE2	8	0	DC	0V
*
* MOTOR POSITION
FPOS	0	11	VSENSE2	1
CPOS	11	0	1
RPOS	11	0	1MEG
*
* ANALYSIS
.TRAN	10MS	200MS
*
* VIEW RESULTS
.PRINT TRAN V(1) I(VSENSE1)
.PROBE
.END
